module Adder1(input [7:0] Ent,
					output[7:0] Sai);			
	assign Sai = Ent + 1'b1;
endmodule