module Instr_Mem( input [7:0]A,
									output reg[31:0]RD);

	always@(*)
	begin
		case(A)
			7'b00000000: 
				RD = 32'b001000_00000_00001_0000000000000011;
			7'b00000001: 
				RD = 32'b00100000000000100000000000001001;
			7'b00000010: 
				RD = 32'b00000000001000100001000000100000;
			7'b00000011: 
				RD = 32'b00000000001000100001100000100100;
			7'b00000100: 
				RD = 32'b00000000001000100010000000100101;
			7'b00000101: 
				RD = 32'b00000000001000100011000000101010;
			7'b00000110: 
				RD = 32'b00000000010000010011100000101010;
			default: 
				RD = 32'b00000000000000000000000000000000;
		endcase
	end

endmodule
